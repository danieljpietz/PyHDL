{name}: if {condition} then
{if_str}
{else_str}
end if {name};