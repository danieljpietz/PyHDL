package {name} is
{types}
{constants}
{procedures}
end package {name};