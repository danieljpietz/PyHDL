function {name} ({args}) return {ret_type} is
begin
{body}
end {name};