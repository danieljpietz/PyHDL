entity {name} is
	port ({interfaces});
end entity {name};