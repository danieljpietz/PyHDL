procedure {name} ({interfaces}) is
{declarations}
begin
{body}
end procedure {name};