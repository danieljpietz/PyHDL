if {condition} then
{body}
end if;