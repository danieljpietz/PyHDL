entity {name} is
end entity {name};