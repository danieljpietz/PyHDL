architecture {name} of {entity} is
{declarations}
begin
{functionality}
end architecture {name};