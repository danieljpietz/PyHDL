component {name} is
	port ({interfaces});
end component {name};