{name}: if {condition} then
{body}
end if {name};