{name} : process {sensitivity}
begin
{body}
end process {name};