package {name} is
{types}
{constants}
end package {name};